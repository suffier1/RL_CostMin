module top_1598227639_809568180_776209382_1234615 (a, b, c, d, e, f, g, h, o);
 input a, b, c, d, e, f, g, h;
 output o;
 and_1 g0(a,b,y1);
 and_1 g1(1'b0,y1,y2);
 and_1 g2(d,y2,y3);
 and_1 g3(e,y3,y4);
 and_1 g4(f,y4,y5);
 and_1 g5(g,y5,y6);
 and_1 g6(h,y6,o);
endmodule
