module top_1598227639_809568180_776209382_1234615 (a, b, c, d, e, f, g, h, o);
 input a, b, c, d, e, f, g, h;
 output o;
 and_1 g0(a,b,y1);
 and_1 g1(1'b0,d,y2);
 and_1 g2(e,f,y3);
 and_1 g3(g,h,y4);
 and_1 g4(y1,y2,y5);
 and_1 g5(y3,y4,y6);
 and_1 g6(y5,y6,o);
endmodule
